`timescale 1ns / 1ps
// `define PRETRAINED

module testbench ( );

	parameter CLOCK_PERIOD = 10;

	logic CLOCK_50;
    logic [0:0] KEY;
    logic [6:0] HEX0;

	// Neuron Test
	logic 				reset;
	logic [15:0] 		neuronIn;
	logic [15:0] 		neuronOut;
	logic 				neuronValid;
	logic 				neuronOutValid;

    // Serializer Test
    parameter numInputs = 784;
    parameter dataWidth = 16;
    parameter counterWidth = $clog2(numInputs);
    logic [numInputs*dataWidth-1:0] inputData;
    logic [dataWidth-1:0] serializerOut;
    logic [counterWidth-1:0] counterOut;
    logic counterValid;


    // Weight Memory
    logic [15:0]       weightMem [0:numInputs-1];

    initial begin
        $readmemb("weight_L0_N0.mif", weightMem);
        $display("Loaded weights:");
        for (int i = 0; i < 16; i++)
            $display("weightMem[%0d] = %b", i, weightMem[i]);
    end

	initial begin
        CLOCK_50 <= 1'b0;
	end // initial
	always @ (*)
	begin : Clock_Generator
		#((CLOCK_PERIOD) / 2) CLOCK_50 <= ~CLOCK_50;
	end
	
	initial begin
        reset <= 1'b0;
        #10
        reset <= 1'b1;
		#10 
		reset <= 1'b0;
		inputData <= 'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000015102e7027e025e00f100910000000000000000000000000000000000000000000000000000000000000000000000000000000000000000037b03fc03fc03fc03fc03c8031b031b031b031b031b031b031b031b02ab00d1000000000000000000000000000000000000000000000000010d01ca012101ca028f039003fc038803fc03fc03fc03ec039803fc03fc023200000000000000000000000000000000000000000000000000000000000000000000004401090038010d010d010d00ed005403b403fc01aa000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000014d03f80347004800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000005803a80400014d000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020603fc03bc00b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ed03e803fc00f9000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000021603fc02ef0014000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000024033703e400e900000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001fa03fc02db000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000012d03f003c400e500000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c037703fc029b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c032f03fc036f008d00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000009903fc03fc013500000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007c038403fc01ce000400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000021603fc03fc00d10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000f503cc03fc03fc00d10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001e603fc03fc036f00a10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001e603fc033f0048000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
        ;   
        #20
		neuronValid <= 1'b1;
        
	end // initial

    always_ff @(posedge CLOCK_50) begin
        if (neuronOutValid)
            $display("Time=%t | neuronOut = %h", $time, neuronOut);
    end

	
	neuron #(
        .layerNumber(0),
        .neuronNumber(0),
        .numWeights(numInputs),
        .dataWidth(dataWidth),
        .dataIntWidth(8),
        .dataFracWidth(8),
        .weightWidth(16),
        .weightIntWidth(8),
        .weightFracWidth(8),
        .biasFile("bias_L0_N0.mif"),
        .weightFile("weight_L0_N0.mif")
    ) U1 (
        .clk(CLOCK_50),
        .reset(reset),
        .neuronIn(serializerOut),
        .neuronValid(neuronValid),
        .weightValid(),
        .weightWriteEn(),
        .biasWriteEn(),
        .weightData(32'h0),
        .biasData(32'h0),
        .config_layer_number(32'h0),
        .config_neuron_number(32'h0),
        .neuronOut(neuronOut),
        .neuronOutValid(neuronOutValid)
    );

     // Serializer Instance
    inputSerializer #(
        .numInputs(numInputs), 
        .dataWidth(dataWidth), 
        .counterWidth(counterWidth)
    ) serializer (
        .clk(CLOCK_50),
        .reset(reset),
        .enable(neuronValid),
        .serializerIn(inputData),
        .counterValid(counterValid),
        .serializerOut(serializerOut)
    );

endmodule
