module NeuralNetwork #(
    parameter   numInputs = 784, numOutputs = 10, L0neurons = 16, L1neurons = 10,
                dataWidth = 16, dataIntWidth = 8, dataFracWidth = 8,
                weightWidth = 16, weightIntWidth = 8, weightFracWidth = 8
) (
    input   logic                               clk,
    input   logic                               reset, 
    input   logic   [dataWidth*numInputs-1:0]   NNin,
    input   logic                               NNvalid,

    output  logic   [dataWidth*numOutputs-1:0]  NNout,
    output  logic                               NNoutValid,
    output  logic   [3:0]                       maxIndex,
    output  logic   [dataWidth-1:0]             maxValue,
    output  logic                               maxValid

);

logic [dataWidth*L0neurons-1:0] layer0Out;
logic                           layer0OutValid;
logic [dataWidth*L1neurons-1:0] layer1Out;
logic                           layer1OutValid;

// logic   [dataWidth*numInputs-1:0]   NNinTest;

// assign NNinTest = 'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000A8B173713F412F30788048500000000000000000000000000000000000000000000000000000000000000000000000000000000000000001BDC1FE01FE01FE01FE01E3E18D918D918D918D918D918D918D918D91555068700000000000000000000000000000000000000000000000008680E4E09090E4E14741C7C1FE01C3C1FE01FE01FE01F5F1CBD1FE01FE01192000000000000000000000000000000000000000000000000000000000000000000000222084801C2086808680868076702A31D9E1FE00D4D0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000A6A1FC01A3A02420000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002C31D3D20000A6A00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010301FE01DDE05860000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007671F3F1FE007C800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010B11FE0177700A100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000012119BA1F1F07470000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FD01FE016D700000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000009691F7F1E1E07270000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002621BBC1FE014D500000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000006019791FE01B7B04640000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004C51FE01FE009AA0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003E41C1C1FE00E6E00200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010B11FE01FE006870000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007A81E5E1FE01FE00687000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000F2F1FE01FE01B7B0505000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000F2F1FE019FA0242000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// assign NNinTest = 'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000100010001000100010001000100010001000100010000000000000000000000000000000000000000000000000000000000000000000000010001000100010001000100010001000100010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;


layer0 #(
    .layerNumber(0), 
    .numInputs(numInputs), 
    .numNeurons(L0neurons),
    .dataWidth(dataWidth), 
    .dataIntWidth(dataIntWidth),
    .dataFracWidth(dataFracWidth),
    .weightWidth(weightWidth),
    .weightIntWidth(weightIntWidth),
    .weightFracWidth(weightFracWidth)
) layer0_inst (
    // Inputs
    .clk(clk),
    .reset(reset),
    .layerIn(NNin),
    .layerValid(NNvalid),
    // Outputs
    .layerOut(layer0Out),
    .layerOutValid(layer0OutValid)
);

layer1 #(
    .layerNumber(1), 
    .numInputs(L0neurons), 
    .numNeurons(L1neurons),
    .dataWidth(dataWidth), 
    .dataIntWidth(dataIntWidth),
    .dataFracWidth(dataFracWidth),
    .weightWidth(weightWidth),
    .weightIntWidth(weightIntWidth),
    .weightFracWidth(weightFracWidth)
) layer1_inst (
    // Inputs
    .clk(clk),
    .reset(reset),
    .layerIn(layer0Out),
    .layerValid(layer0OutValid),
    // Outputs
    .layerOut(NNout),
    .layerOutValid(NNoutValid)
);

hardmax #(
    .dataWidth(dataWidth), 
    .numOutputs(10)
) hardmax_inst (
    // Inputs
    .clk(clk),
    .reset(reset),
    .dataIn(NNout),
    .enable(NNoutValid),
    // Outputs
    .maxIndex(maxIndex),
    .maxValue(maxValue),
    .maxValid(maxValid)
);
    
endmodule