`timescale 1ns / 1ps
// `define PRETRAINED

module testbench ( );

	parameter CLOCK_PERIOD = 10;

	logic CLOCK_50;
    logic [0:0] KEY;
    logic [6:0] HEX0;

	// Neuron Test
	logic 				reset;
	logic [15:0] 		neuronIn;
	logic [15:0] 		neuronOut;
	logic 				neuronValid;
	logic 				neuronOutValid;

    // Serializer Test
    parameter numInputs = 784;
    parameter dataWidth = 16;
    parameter counterWidth = $clog2(numInputs);
    logic [numInputs*dataWidth-1:0] inputData;
    logic [dataWidth-1:0] serializerOut;
    logic [counterWidth-1:0] counterOut;
    logic counterValid;


    // Weight Memory
    logic [15:0]       weightMem [0:numInputs-1];

    initial begin
        $readmemb("weight_L0_N0.mif", weightMem);
        $display("Loaded weights:");
        for (int i = 0; i < 16; i++)
            $display("weightMem[%0d] = %b", i, weightMem[i]);
    end

	initial begin
        CLOCK_50 <= 1'b0;
	end // initial
	always @ (*)
	begin : Clock_Generator
		#((CLOCK_PERIOD) / 2) CLOCK_50 <= ~CLOCK_50;
	end
	
	initial begin
        reset <= 1'b0;
        #10
        reset <= 1'b1;
		#10 
		reset <= 1'b0;
		inputData <= 'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000A8B173713F412F30788048500000000000000000000000000000000000000000000000000000000000000000000000000000000000000001BDC1FE01FE01FE01FE01E3E18D918D918D918D918D918D918D918D91555068700000000000000000000000000000000000000000000000008680E4E09090E4E14741C7C1FE01C3C1FE01FE01FE01F5F1CBD1FE01FE01192000000000000000000000000000000000000000000000000000000000000000000000222084801C2086808680868076702A31D9E1FE00D4D0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000A6A1FC01A3A02420000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002C31D3D20000A6A00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010301FE01DDE05860000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007671F3F1FE007C800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010B11FE0177700A100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000012119BA1F1F07470000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FD01FE016D700000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000009691F7F1E1E07270000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002621BBC1FE014D500000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000006019791FE01B7B04640000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004C51FE01FE009AA0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003E41C1C1FE00E6E00200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010B11FE01FE006870000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007A81E5E1FE01FE00687000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000F2F1FE01FE01B7B0505000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000F2F1FE019FA0242000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
        ;
        #20
		neuronValid <= 1'b1;
        
	end // initial

    always_ff @(posedge CLOCK_50) begin
        if (neuronOutValid)
            $display("Time=%t | neuronOut = %h", $time, neuronOut);
    end

	
	neuron #(
        .layerNumber(0),
        .neuronNumber(0),
        .numWeights(numInputs),
        .dataWidth(dataWidth),
        .dataIntWidth(8),
        .dataFracWidth(8),
        .weightWidth(16),
        .weightIntWidth(8),
        .weightFracWidth(8),
        .biasFile("bias_L0_N0.mif"),
        .weightFile("weight_L0_N0.mif")
    ) U1 (
        .clk(CLOCK_50),
        .reset(reset),
        .neuronIn(serializerOut),
        .neuronValid(neuronValid),
        .weightValid(),
        .weightWriteEn(),
        .biasWriteEn(),
        .weightData(32'h0),
        .biasData(32'h0),
        .config_layer_number(32'h0),
        .config_neuron_number(32'h0),
        .neuronOut(neuronOut),
        .neuronOutValid(neuronOutValid)
    );

     // Serializer Instance
    inputSerializer #(
        .numInputs(numInputs), 
        .dataWidth(dataWidth), 
        .counterWidth(counterWidth)
    ) serializer (
        .clk(CLOCK_50),
        .reset(reset),
        .enable(neuronValid),
        .serializerIn(inputData),
        .counterValid(counterValid),
        .serializerOut(serializerOut)
    );

endmodule
