`timescale 1ns / 1ps
// `define PRETRAINED

module testbench ( );

	parameter CLOCK_PERIOD = 10;
    parameter NUM_INPUTS = 784;
    parameter NUM_NEURONS = 16;
    parameter DATA_WIDTH = 16;

	logic CLOCK_50;

	// Layer Test
	logic 				reset;
	logic [NUM_INPUTS*DATA_WIDTH-1:0] 		layerIn;
	logic [NUM_NEURONS*DATA_WIDTH-1:0] 		layerOut;
	logic 				layerValid;
	logic 				layerOutValid;

    // Weight Memory
    logic [DATA_WIDTH-1:0]       weightMem [0:255];


    initial begin
        $readmemb("weights/weight_L0_N0.mif", weightMem);
        $display("Loaded weights:");
        for (int i = 0; i < 16; i++)
            $display("weightMem[%0d] = %b", i, weightMem[i]);
    end

	initial begin
        CLOCK_50 <= 1'b0;
	end // initial
	always @ (*)
	begin : Clock_Generator
		#((CLOCK_PERIOD) / 2) CLOCK_50 <= ~CLOCK_50;
	end
	
	initial begin
        reset <= 1'b0;
        // layerIn <= {392{16'h0203}};
        //'h297F3C12A49D562B00FF1A4E9063C1887634204599AFBE1867D32C4AE207851E543DA8910CF2B46B1D7E39C7E14028ABFC0F3E5D2A8473656E89A210B5374F9B0B112233445566778899AABBCCDDEEFFFEDCBA98765432100123456789ABCDEFC0C1C2C3C4C5C6C7C8C9CACBCCCDCECFD0D1D2D3D4D5D6D7D8D9DADBDCDDDEDFE0E1E2E3E4E5E6E7E8E9EAEBECEDEEF0F1F2F3F4F5F6F7F8F9FAFBFCFDFEFF000102030405060708090A0B0C0D0E0F101112131415161718191A1B1C1D1E1F202122232425262728292A2B2C2D2E2F303132333435363738393A3B3C3D3E3F404142434445464748494A4B4C4D4E4F505152535455565758595A5B5C5D5E5F606162636465666768696A6B6C6D6E6F707172737475767778797A7B7C7D7E7F808182838485868788898A8B8C8D8E8F909192939495969798999A9B9C9D9E9FA0A1A2A3A4A5A6A7A8A9AAABACADAEAFB;
        layerIn <= 'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000015102e7027e025e00f100910000000000000000000000000000000000000000000000000000000000000000000000000000000000000000037b03fc03fc03fc03fc03c8031b031b031b031b031b031b031b031b02ab00d1000000000000000000000000000000000000000000000000010d01ca012101ca028f039003fc038803fc03fc03fc03ec039803fc03fc023200000000000000000000000000000000000000000000000000000000000000000000004401090038010d010d010d00ed005403b403fc01aa000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000014d03f80347004800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000005803a80400014d000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020603fc03bc00b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ed03e803fc00f9000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000021603fc02ef0014000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000024033703e400e900000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001fa03fc02db000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000012d03f003c400e500000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c037703fc029b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c032f03fc036f008d00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000009903fc03fc013500000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007c038403fc01ce000400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000021603fc03fc00d10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000f503cc03fc03fc00d10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001e603fc03fc036f00a10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001e603fc033f0048000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
        ;
        #10
        reset <= 1'b1;
		#10 
		reset <= 1'b0;
		#10
		layerValid <= 1'b1;
	end // initial

    layer #(
        .layerNumber(0),
        
        .numInputs(NUM_INPUTS),
        .numNeurons(NUM_NEURONS),
        .dataWidth(DATA_WIDTH),
        .dataIntWidth(6),
        .dataFracWidth(10),
        .weightWidth(DATA_WIDTH),
        .weightIntWidth(6),
        .weightFracWidth(10)

    ) U1 (
        .clk(CLOCK_50),
        .reset(reset),
        .layerIn(layerIn),
        .layerValid(layerValid),
        .layerOut(layerOut),
        .layerOutValid(layerOutValid)
    );

endmodule
