`timescale 1ns / 1ps
// `define PRETRAINED

module testbench ( );

	parameter CLOCK_PERIOD = 10;
    parameter SCLK = 15;

	// top Test
	logic 				reset;
	logic               CLOCK_50;
    logic               serialClock;
    logic               serialData;
    logic   [6:0]       HEX0;
    logic   [1:0]       KEY;
    logic   [15:0]      ARDUINO_IO;


    logic   [784*16-1:0]    data;

	initial begin
        CLOCK_50 <= 1'b0;
        serialClock <= 1'b0;
	end // initial
	always @ (*)
	begin : Clock_Generator
		#((CLOCK_PERIOD) / 2) CLOCK_50 <= ~CLOCK_50;
	end
    always @ (*)
	begin : Clock_Generator_2
		#((SCLK) / 2) serialClock <= ~serialClock;
	end

    integer i;
	
	initial begin
        data = 'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000A8B173713F412F30788048500000000000000000000000000000000000000000000000000000000000000000000000000000000000000001BDC1FE01FE01FE01FE01E3E18D918D918D918D918D918D918D918D91555068700000000000000000000000000000000000000000000000008680E4E09090E4E14741C7C1FE01C3C1FE01FE01FE01F5F1CBD1FE01FE01192000000000000000000000000000000000000000000000000000000000000000000000222084801C2086808680868076702A31D9E1FE00D4D0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000A6A1FC01A3A02420000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002C31D3D20000A6A00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010301FE01DDE05860000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007671F3F1FE007C800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010B11FE0177700A100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000012119BA1F1F07470000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FD01FE016D700000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000009691F7F1E1E07270000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002621BBC1FE014D500000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000006019791FE01B7B04640000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004C51FE01FE009AA0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003E41C1C1FE00E6E00200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010B11FE01FE006870000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007A81E5E1FE01FE00687000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000F2F1FE01FE01B7B0505000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000F2F1FE019FA0242000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        reset <= 1'b0;
        #10
        reset <= 1'b1;
		#10 
		reset <= 1'b0;
		#10
		for (i = 0; i < 784 * 16; i = i + 1) begin
            serialData <= data[i];
            #15;
        end
	end // initial

    top U1 (
        .KEY({~reset,1'b0}),
        .CLOCK_50(CLOCK_50),
        .HEX0(HEX0),
        .ARDUINO_IO({14'b0, serialData, serialClock})
    ); 

endmodule
