`timescale 1ns / 1ps
// `define PRETRAINED

module testbench ( );

	parameter CLOCK_PERIOD = 10;

	logic CLOCK_50;

	// Layer Test
	logic 				reset;
	logic [784*8-1:0] 	NNin;
	logic [10*8-1:0] 	NNout;
	logic 			    NNvalid;
	logic 			    NNoutValid;
    logic [3:0]         maxIndex;
    logic [7:0]         maxValue;
    logic               maxValid;

    // Memory
    logic [784*8-1:0] mem [0:7];
    initial begin
        $readmemh("flattened_inputs_hex.mif", mem);
    end

	initial begin
        CLOCK_50 <= 1'b0;
	end // initial
	always @ (*)
	begin : Clock_Generator
		#((CLOCK_PERIOD) / 2) CLOCK_50 <= ~CLOCK_50;
	end
	
	initial begin
        reset <= 1'b0;
        //NNin <= 6272'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002a5d504c1e12000000000000000000000000000000000000000000006f7f7f7f7f796363636363636363551a0000000000000000000000002239243952727f717f7f7f7d737f7f4600000000000000000000000000000000000921072222221e0b767f350000000000000000000000000000000000000000000000002a7f690900000000000000000000000000000000000000000000000b757f2a000000000000000000000000000000000000000000000000417f771600000000000000000000000000000000000000000000001e7d7f1f000000000000000000000000000000000000000000000000437f5e03000000000000000000000000000000000000000000000005677c1d0000000000000000000000000000000000000000000000003f7f5b000000000000000000000000000000000000000000000000267e781d00000000000000000000000000000000000000000000000a6f7f53000000000000000000000000000000000000000000000002667f6e120000000000000000000000000000000000000000000000137f7f27000000000000000000000000000000000000000000000010707f3a010000000000000000000000000000000000000000000000437f7f1a00000000000000000000000000000000000000000000001f797f7f1a00000000000000000000000000000000000000000000003d7f7f6e1400000000000000000000000000000000000000000000003d7f6809000000000000000000000000000000000000000000000000000000000000000000000000000000000000
        //NNin <= 6272'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003a3f567f7f4b2f0000000000000000000000000000000000000000557f7f7f7f7f7f6d0f000000000000000000000000000000000000557f7f7f6b47587f7f3d00000000000000000000000000000000001a7d7f6910060003677f460000000000000000000000000000000000277e690d0000003d7c7f21000000000000000000000000000000000000100900000000697f7f2100000000000000000000000000000000000000000000003b7c7f630500000000000000000000000000000000000000000000267c7f74200000000000000000000000000000000000000000000000407f7f480000000000000000000000000000000000000000000000587b7f5006000000000000000000000000000000000000000000000d757f75120000000000000000000000000000000000000000000000637f7f470000000000000000000000000000000000000000000000277c7f5f06000000000000000000000000000000000000000000000a647f7f470000000000000000000000000000000000000000000000437f7f570600000000000000000000000000000000000000000000007c7f7f0d0000000000000000000000000000000000000000000000007c7f7f160a0a0a0a0300030a0a134b4b4b4a050000000000000000007c7f7f7f7f7f7f7f5448537f7f7f7f7f7f7f3e000000000000000000577f7f7f7f7f7f7f7f7f7f7f7d7c7c553b3b1d000000000000000000003b3e3e3e537f7f7f4e3e3e15000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
        //NNin <= 6272'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000137f37000000000000000000000000000000000000000000000000002c7e2900000000000000000000000000000000000000000000000000447900000000000000000000000000000000000000000000000000177a4b000000000000000000000000000000000000000000000000002a7f2000000000000000000000000000000000000000000000000000657006000000000000000000000000000000000000000000000000107f6c00000000000000000000000000000000000000000000000000307f6200000000000000000000000000000000000000000000000000467f270000000000000000000000000000000000000000000000001d7767040000000000000000000000000000000000000000000000003e7f5300000000000000000000000000000000000000000000000000567f290000000000000000000000000000000000000000000000000c746c000000000000000000000000000000000000000000000000003c7f50000000000000000000000000000000000000000000000000004c7f4700000000000000000000000000000000000000000000000000727f210000000000000000000000000000000000000000000000001f7e7f21000000000000000000000000000000000000000000000000477f67020000000000000000000000000000000000000000000000056c7f3d00000000000000000000000000000000000000000000000003635805000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
        //NNin <= 6272'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000064b7f65100000000000000000000000000000000000000000000000137e7e7f36000000000000000000000000000000000000000000000b637e7e7f36000000000000000000000000000000000000000000375f7e7e7e7f55371f000000000000000000000000000000000000007f7e7e7e7e7f7e7e6e1a00000000000000000000000000000000005b7f7f7f7f7f756f7f7f7f00000000000000000000000000000000206f7f7e7e7e4a271f407e7e35000000000000000000000000000010747e7f7e6e4505000010737e7a3903000000000000000000000000137e7e7f5e0a0000000000377e7f7e12000000000000000000000000137e7e650f00000000000010647f7e12000000000000000000000000137f7f000000000000000010657f7f52000000000000000000000000467e7e0000000000000000377e7f7e120000000000000000000000006d7e7e0000000000000b20747e7f730f0000000000000000000000006d7e7e000000000000487e7e7e6f1f000000000000000000000000006d7e7e00000000005b6f7e7e7e5a00000000000000000000000000006d7f7f2525727f7f7f7f7f7f7f000000000000000000000000000000397e7e7f7e7e7e7e7f7e7e7e4a00000000000000000000000000000010737e7f7e7e7e7e7f735f1205000000000000000000000000000000001f477f7e7e7e7e7f3600000000000000000000000000000000000000000024577e5724240f000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
        //NNin <= 6272'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000074b610300000000000000000000000000000000000000000000002e707f7f0a000000000000000000000000000000000000000000000e767f7f7f5309000000000000000000000000000000000000000000487f7f7f7f7f773a0300000000000000000000000000000000000010797f685d7f7f7f740c000000000000000000000000000000000000287f610004316e7f7f650900000000000000000000000000000000002b7f280000005b7f7f60060000000000000000000000000000000000587f4e000000757f7f440000000000000000000000000000000000002b7f68142b537e777f7615000000000000000000000000000000000009777f7f7f7f5d126c7f4c00000000000000000000000000000000000022787f7f490400437f7012000000000000000000000000000000000000224f4706000005587f51000000000000000000000000000000000000000000000000002c7f710900000000000000000000000000000000000000000000000001537f3f00000000000000000000000000000000000000000000000000187b7f13000000000000000000000000000000000000000000000000003a7f56050000000000000000000000000000000000000000000000000b6d7f17000000000000000000000000000000000000000000000000000f7f5300000000000000000000000000000000000000000000000000005d7a1500000000000000000000000000000000000000000000000000077027000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
        //NNin <= 6272'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000b604310000000000000000008270300000000000000000000000009767d550000000000000000086e791300000000000000000000000a5f7f4a000000000000000000467f32000000000000000000000000237f7f0b0000000000000000167f570700000000000000000000000b4d7f30000000000000000016747f2e000000000000000000000000527f66060000000000000000347f4f00000000000000000000000000517f59030000000000000542777f0000000000000000000000000000517f7f60582323232343637f7f5500000000000000000000000000001a727f7f7f7f7f7f7f7f7f7f6e120000000000000000000000000000000921457f74454545167f7f51000000000000000000000000000000000000000000000000117f670b000000000000000000000000000000000000000000000000507f230000000000000000000000000000000000000000000000002b7f79190000000000000000000000000000000000000000000000004f7f5300000000000000000000000000000000000000000000000000747a19000000000000000000000000000000000000000000000000347f7400000000000000000000000000000000000000000000000000687f4f00070f00000000000000000000000000000000000000000000687f4d2e665100000000000000000000000000000000000000000000687f7f7f4d0f000000000000000000000000000000000000000000001f5f400c0300000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
        NNin <= mem[1]; // Load the first input from memory
        #10
        reset <= 1'b1;
		#10 
		reset <= 1'b0;
		#10
		NNvalid <= 1'b1;
	end // initial

    NeuralNetwork #(
        .dataWidth(8), 
        .numInputs(784), 
        .numOutputs(10), 
        .L0neurons(16), 
        .L1neurons(10)
    ) nn (
        .clk(CLOCK_50),
        .reset(reset),
        .NNin(NNin),
        .NNvalid(NNvalid),
        .NNout(NNout),
        .NNoutValid(NNoutValid),
        .maxIndex(maxIndex),
        .maxValid(maxValid),
        .maxValue(maxValue)
    );

endmodule
